entity deneme is
end entity;

architecture sim of deneme is
begin

    process is 
    begin
        report "Hello World";
        wait;

    end process;

end architecture;